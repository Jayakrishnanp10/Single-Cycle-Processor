module instruction_memory( input [31:0]A,
		output reg [31:0]RD);

reg [7:0] REG [65535:0];

always @(A) begin
RD<={REG[A+32'h00000003],REG[A+32'h00000002],REG[A+32'h00000001],REG[A]};
	    
end

assign {REG[32'h00001003],REG[32'h00001002],REG[32'h00001001],REG[32'h00001000]} = 32'hFFC4A303;
assign {REG[32'h00001007],REG[32'h00001006],REG[32'h00001005],REG[32'h00001004]} = 32'h0064A423;
assign {REG[32'h0000100B],REG[32'h0000100A],REG[32'h00001009],REG[32'h00001008]} = 32'h0062E233;
assign {REG[32'h0000100F],REG[32'h0000100E],REG[32'h0000100D],REG[32'h0000100C]} = 32'hFDA48393;
assign {REG[32'h00001013],REG[32'h00001012],REG[32'h00001011],REG[32'h00001010]} = 32'hFE420AE3;
endmodule

